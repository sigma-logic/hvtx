// Copyright (c) 2025 Sigma Logic

`include "h14tx/registers.svh"

// Implementation of HDMI Auxiliary Video InfoFrame packet.
// By Sameer Puri https://github.com/sameer

// See Section 8.2.1
module h14tx_pkt_avi_info_frame
    import h14tx_pkg::packet_t;
#(
    parameter bit [1:0] VideoFormat = 2'b00,  // 00 = RGB, 01 = YCbCr 4:2:2, 10 = YCbCr 4:4:4
    parameter bit ActiveFormatInfoPresent = 1'b0,  // Not valid
    parameter bit [1:0] BarInfo = 2'b00,  // Not valid
    parameter bit [1:0] ScanInfo = 2'b00,  // No data
    parameter bit [1:0] Colorometry = 2'b00,  // No data
    parameter bit [1:0] PictureAspectRatio = 2'b00, // No data, See CEA-CEB16 for more information about Active Format Description processing.
    parameter bit [3:0] ActiveFormatAspectRatio = 4'b1000, // Not valid unless ActiveFormatInfoPresent = 1'b1, then Same as picture aspect ratio
    parameter bit ItContent = 1'b0, //  The IT content bit indicates when picture content is composed according to common IT practice (i.e. without regard to Nyquist criterion) and is unsuitable for analog reconstruction or filtering. When the IT content bit is set to 1, downstream processors should pass pixel data unfiltered and without analog reconstruction.
    parameter bit [2:0] ExtendedColorometry = 3'b000, // Not valid unless Colorometry = 2'b11. The extended colorimetry bits, EC2, EC1, and EC0, describe optional colorimetry encoding that may be applicable to some implementations and are always present, whether their information is valid or not (see CEA 861-D Section 7.5.5).
    parameter bit [1:0] RgbQuantizationRange = 2'b00, // Default. Displays conforming to CEA-861-D accept both a limited quantization range of 220 levels (16 to 235) anda full range of 256 levels (0 to 255) when receiving video with RGB color space (see CEA 861-D Sections 5.1, Section 5.2, Section 5.3 and Section 5.4). By default, RGB pixel data values should be assumed to have the limited range when receiving a CE video format, and the full range when receiving an IT format. The quantization bits allow the source to override this default and to explicitly indicate the current RGB quantization range.
    parameter bit [1:0] NonUniformPictureScaling = 2'b00, // None. The Nonuniform Picture Scaling bits shall be set if the source device scales the picture or has determined that scaling has been performed in a specific direction.
    parameter int VideoIdCode = 4,  // Same as the one from the HDMI module
    parameter bit [1:0] YccQuantizationRange = 2'b00,  // 00 = Limited, 01 = Full
    parameter bit [1:0] ContentType = 2'b00,  // No data, becomes Graphics if ItContent = 1'b1.
    parameter bit [3:0] PixelRepetition = 4'b0000  // None
) (
    output packet_t packet
);

    localparam bit [4:0] Length = 5'd13;
    localparam bit [7:0] Version = 8'd2;
    localparam bit [6:0] Type = 7'd2;

    assign packet.header = {{3'b0, Length}, Version, {1'b1, Type}};

    // PB0-PB6 = sub0
    // PB7-13 =  sub1sus
    // PB14-20 = sub2
    // PB21-27 = sub3
    logic [7:0] packet_bytes[27:0];

    assign packet_bytes[0] = 8'd1 + ~(packet.header[23:16] + packet.header[15:8] + packet.header[7:0] + packet_bytes[13] + packet_bytes[12] + packet_bytes[11] + packet_bytes[10] + packet_bytes[9] + packet_bytes[8] + packet_bytes[7] + packet_bytes[6] + packet_bytes[5] + packet_bytes[4] + packet_bytes[3] + packet_bytes[2] + packet_bytes[1]);
    assign packet_bytes[1] = {1'b0, VideoFormat, ActiveFormatInfoPresent, BarInfo, ScanInfo};
    assign packet_bytes[2] = {Colorometry, PictureAspectRatio, ActiveFormatAspectRatio};
    assign packet_bytes[3] = {
        ItContent, ExtendedColorometry, RgbQuantizationRange, NonUniformPictureScaling
    };
    assign packet_bytes[4] = {1'b0, 7'(VideoIdCode)};
    assign packet_bytes[5] = {YccQuantizationRange, ContentType, PixelRepetition};

    genvar i;
    generate
        // Assign values to bars if BAR_INFO says they are valid
        if (BarInfo != 2'b00) begin
            assign packet_bytes[6]  = 8'hff;
            assign packet_bytes[7]  = 8'hff;
            assign packet_bytes[8]  = 8'h00;
            assign packet_bytes[9]  = 8'h00;
            assign packet_bytes[10] = 8'hff;
            assign packet_bytes[11] = 8'hff;
            assign packet_bytes[12] = 8'h00;
            assign packet_bytes[13] = 8'h00;
        end else begin
            assign packet_bytes[6]  = 8'h00;
            assign packet_bytes[7]  = 8'h00;
            assign packet_bytes[8]  = 8'h00;
            assign packet_bytes[9]  = 8'h00;
            assign packet_bytes[10] = 8'h00;
            assign packet_bytes[11] = 8'h00;
            assign packet_bytes[12] = 8'h00;
            assign packet_bytes[13] = 8'h00;
        end
        for (i = 14; i < 28; i++) begin : pb_reserved
            assign packet_bytes[i] = 8'd0;
        end
        for (i = 0; i < 4; i++) begin : pb_to_sub
            assign packet.sub[i] = {
                packet_bytes[6+i*7],
                packet_bytes[5+i*7],
                packet_bytes[4+i*7],
                packet_bytes[3+i*7],
                packet_bytes[2+i*7],
                packet_bytes[1+i*7],
                packet_bytes[0+i*7]
            };
        end
    endgenerate

endmodule

