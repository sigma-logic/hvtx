module dev();
endmodule : dev
