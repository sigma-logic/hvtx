`ifndef H14TX_TYPEDEFS_SVH_
`define H14TX_TYPEDEFS_SVH_

`endif
