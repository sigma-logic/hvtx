`ifndef H14TX_MACROS_SVH_
`define H14TX_MACROS_SVH_

`define VEC(width) logic [width-1:0]

`endif
